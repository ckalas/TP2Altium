*****************************************************************
* SPICE2G6 MODEL OF THE DIODE BAW101  (SOT-23)                  *
* REV: 98.1                  DANALYSE GMBH BERLIN (27.07.1998)  *
*****************************************************************
* jjt 31/10/2000: moved the model into the subckt
*
.SUBCKT BAW101 1 2
D    3 4 DBAW101
L1   1 3 0.350N
L2   4 2 0.350N
.MODEL DBAW101 D
+ IS  =  0.2583E-12
+ N   =  1.1790
+ RS  =  3.0000
+ EG  =  1.1073
+ XTI =  4.4349
+ CJO =  6.2000E-12
+ VJ  =  0.7000
+ M   =  0.5000
.ENDS
