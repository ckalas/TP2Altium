*****************************************************************
.SUBCKT BAT17-05W 1 2 3
D1 1 3 D188
D2 2 3 D188
.MODEL D188 D(IS=4n RS=3.3 N=1.03 XTI=2 EG=.65
+ CJO=415f M=.156 VJ=.115 FC=.5 BV=12 IBV=5U TT=25p)
.ENDS
