*****************************************************************
.SUBCKT BAT68-05 1 2 3
D1 1 3 BAT68
D2 2 3 BAT68
.MODEL BAT68 D(IS=8N RS=2 N=1.05 XTI=1.8 EG=.68
+ CJO=.77P M=.075 VJ=.1 FC=.5 BV=8 IBV=1U TT=25P)
.ENDS
