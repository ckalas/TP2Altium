*****************************************************************
.SUBCKT BAT18-06 1 2 3
D1 3 1 BAT18	
D2 3 2 BAT18
.MODEL BAT18 D(IS=185F RS=.30 N=1.305 BV=70 IBV=.1N
+ CJO=1.17P VJ=.12 M=.096 TT=125N)
.ENDS