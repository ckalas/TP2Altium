*****************************************************************
.SUBCKT BAT66-05 1 2 3
D1 1 2 BAT66
D2 3 2 BAT66
.MODEL BAT66 D(Is=243.5n N=1.001 Rs=0.1401 Xti=3 Eg=1.11 Cjo=170.5p M=0.548
+ Vj=.4803 Fc=.5 Bv=30 Ibv=100u TT=30p)
.ENDS