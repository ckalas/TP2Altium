*****************************************************************
.SUBCKT BAT18-05 1 2 3
D1 1 3 BAT18	
D2 2 3 BAT18
.MODEL BAT18 D(IS=185F RS=.30 N=1.305 BV=70 IBV=.1N
+ CJO=1.17P VJ=.12 M=.096 TT=125N)
.ENDS