******************************************************
.SUBCKT BAV199 1 2 3
D1 1 3 DBAV199
D2 3 2 DBAV199
.MODEL DBAV199 D (IS=510P RS=42M N=1.75 BV=70 IBV=1.4U
+ CJO=2.65P VJ=.75 M=.333 TT=4.32U)
.ENDS BAV199