*****************************************************************
.SUBCKT BAT240A 1 2 3
D1 3 1 D364
D2 1 2 D364
.MODEL D364 D(IS=146N RS=2.18 N=1.07 XTI=4.25 EG=.650 
+ CJO=57.0P M=.495 VJ=.390 FC=.500 BV=240 IBV=5.00U TT=120P)
.ENDS
