***************************************************
.SUBCKT BAR64-06 1 2 3
D1 3 1 BAR64
D2 3 2 BAR64
.MODEL BAR64 D(IS=880p RS=.9 N=1.305 BV=70 IBV=.1N
+ CJO=0.33P VJ=.8 M=.2 TT=1.25u)
.ENDS