*****************************************************************
.SUBCKT BBY52 1 2 3
D1 1 3 D341
D2 2 3 D341
.MODEL D341 D(IS=219E-18 N=1.021 RS=0.4893 XTI=3 EG=1.11 CJO=2.6E-12
+ M=0.452 VJ=0.8 FC=.5 BV=10 IBV=1E-6 TT=120E-9)
.ENDS

* hyperabrupt Diode, M=f(VR)! C-curve approximated between VR=1..6V
* 9.1.96 SIEMENS PD1 Moschovis