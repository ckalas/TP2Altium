*****************************************************************
* SPICE2G6 MODEL OF THE DIODE BAS28W (SOT-23)                    *
* REV: 98.1                  DANALYSE GMBH BERLIN (27.07.1998)  *
*****************************************************************
* jjt 31/10/2000 : moved the model into the subckt
*
.SUBCKT BAS28W 1 2
D    3 4 DBAS28
L1   1 3 0.350N
L2   4 2 0.350N
.MODEL DBAS28 D
+ IS  =  2.7838E-09
+ N   =  1.8703
+ RS  =  1.3548
+ EG  =  1.0637
+ XTI =  1.5000
+ CJO =  0.6000E-12
+ VJ  =  0.2000
+ M   =  0.1000
.ENDS
