*****************************************************************
.SUBCKT BAT15-04W 1 2 3
D1 1 3 BAT15-04
D2 3 2 BAT15-04
.MODEL BAT15-04 D(Is=130n N=1.08 Rs=4.5 Xti=1.8 Eg=.68 Cjo=260f M=.047
+ Vj=.11 Fc=.5 Bv=4 Ibv=10u Tt=25p)
.ENDS

* Case SOT23, 2 diodes, connection pins 1-3 / 3-2
* Data for each diode, add R=3.3MEG parallel to each diode for better IR and
* R0 simulation
* 10.11.1994 SIEMENS HL EH PD1 Kurth