*****************************************************************
.SUBCKT BAS125-04 1 2 3
D1 1 3 BAS125
D2 3 2 BAS125
.MODEL BAS125 D(IS=1.45N RS=12 N=1.03 XTI=1.6 EG=.68
+ CJO=.95P M=.2 VJ=.24 FC=.5 BV=25 IBV=100n TT=25P)
.ENDS

* ISR=15n NR=4k IKF=10m
* for 27C reverse current simulation use GMIN=1e-9

