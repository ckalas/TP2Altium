*****************************************************************
.SUBCKT BAT64-04 1 2 3
D1 1 3 BAT64
D2 3 2 BAT64
.MODEL BAT64 D(
+       AF= 1.00E+00    BV= 3.00E+01   CJO= 6.59E-12    EG= 1.11E+00
+       FC= 5.00E-01   IBV= 1.00E-04    IS= 6.97E-09    KF= 0.00E+00
+        M= 3.96E-01     N= 1.01E+00    RS= 1.84E+00    TT= 1.00E-10
+       VJ= 3.42E-01   XTI= 3.00E+00)
.ENDS