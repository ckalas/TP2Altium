*****************************************************************
.SUBCKT BAR63-06W 1 2 3
D1 3 1 D310
D2 3 2 D310
.model D310 D(Is=60E-18 N=1.02 Rs=.45 Xti=3 Eg=1.11 Cjo=.19p
+ M=.15 Vj=.25 Fc=.5 Bv=50 Ibv=5u Tt=75n)
.ENDS
