*****************************************************************
* SPICE2G6 MODEL OF THE DIODE SMBD7000 (SOT-23)                 *
* REV: 98.1                  DANALYSE GMBH BERLIN (27.07.1998)  *
*****************************************************************
* jjt 31/10/2000: moved model into subckt
*
* Connections:
*                Anode 1
*                | Cathode 2
*                | | Anode 2/Cathode 1
*                | | |
.SUBCKT SMBD7000 1 2 3
X1 1 3 XSMBD7000
X2 3 2 XSMBD7000
.ENDS
.SUBCKT XSMBD7000 1 2
D    3 4 DSMBD7000
L1   1 3 0.350N
L2   4 2 0.350N
.MODEL DSMBD7000 D
+ IS  =  2.7838E-09
+ N   =  1.8703
+ RS  =  1.3548
+ EG  =  1.0637
+ XTI =  1.5000
+ CJO =  0.6000E-12
+ VJ  =  0.2000
+ M   =  0.1000
.ENDS
