*****************************************************************
.SUBCKT BB814 1 2 3
D1 1 3 DBB814
D2 2 3 DBB814
.MODEL DBB814 D(IS=7f N=1.012 RS=.18 XTI=3 EG=1.11 CJO=83.9p M=.775
+ VJ=1.6 FC=.5 BV=20 IBV=100n TT=137n)
.ENDS

*  IKF=1 ISR=10p NR=1K
* hyperabrupt Diode, M=f(VR)! C-curve approximated between VR=1..9V
* BB814-typical, SIEMENS HL EH PD1 KTH 