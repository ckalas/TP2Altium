*****************************************************************
.SUBCKT BAT15-099R 1 2 3 4
D1 1 3 BAT15-099R1
D2 3 2 BAT15-099R1
D3 2 4 BAT15-099R1
D4 4 1 BAT15-099R1
.MODEL BAT15-099R1 D(Is=150n N=1.04 Rs=2.6 Xti=1.8 Eg=.68 Cjo=365f M=.061
+ Vj=.12 Fc=.5 Bv=4 Ibv=10u Tt=25p)
.ENDS

* Case SOT143, 4-diode-chip-ring 1-3-2-4-1, I/O connection 1-2 / 4-3 
* Data for each diode, add R=1.5MEG parallel to each diode for better IR and
* R0 simulation
