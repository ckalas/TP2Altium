*****************************************************************
.SUBCKT BAS40-05W 1 2 3
D1 1 3 BAS40	
D2 2 3 BAS40	
.MODEL BAS40 D(IS=8N RS=7.8 N=1.04 XTI=1.8 EG=.68 
+ CJO=3P M=.42 VJ=.4 FC=.5 BV=40 IBV=100n TT=25P)
.ENDS

* ISR=5n NR=1k IKF=10m
* for 27C reverse current simulation use: GMIN=1e-9
