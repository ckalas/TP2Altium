*****************************************************************
.SUBCKT BBY51 1 2 3
D1 1 3 D340
D2 2 3 D340
.MODEL D340 D(IS=3.3E-15 N=1.115 RS=0.06 XTI=3 EG=1.11 CJO=7.32E-12
+ M=0.914 VJ=2.34 FC=.5 BV=10 IBV=1E-6 TT=5E-9)
.ENDS

* hyperabrupt Diode, M=f(VR)! C-curve approximated between VR=1..6V
* For Capacitance Q-factor add RS=0.44 externally or (degrades VF/IF) 
* internally
* 13.10.95 SIEMENS PD1 KURTH