******************************************************
.SUBCKT BAV170 1 2 3
D1 1 3 DBAV170
D2 2 3 DBAV170
.MODEL DBAV170 D (IS=473P RS=42M N=1.75 BV=70 IBV=1.3U
+ CJO=2.65P VJ=.75 M=.333 TT=4.32U)
.ENDS BAV170
